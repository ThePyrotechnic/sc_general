BZh91AY&SYV�| I߀Py����������`����   U6��2d�@hh@ h ��1D�       9�#� �&���0F&�	�����h2   � 9�#� �&���0F&%4	�114M2��24�f�&��i�ꞓ�?Tв�{D�LT?��)FȒ�%?H!`�"�"�BT+��P܂co">��	�LLeOi�K�l�W����:%Hϴn���إ�RhA���ԁ
�eb��]�[ɺ���:���l�[�L��"t��f�F��!B,��'!�f�\�����n[-��,ӑ� �M��r���0C0����F�Z��B�B~��@u�C$��=����p"x=�P��e�A2�e�ir��d�c�E���d���:����Q���M�l��� Z�ũGL,ӆ�̣55C}��E��C"���������di@���&aUق�V�G�  ���L9�7�&J4Ņ��� ��ZT�I����kDT�ł=h,�t�-I��C�C0�[Af�${"K0E�&���6��T)0d��F��%&�.���9�BBt�$	$H!E�.�iԀ��"����#2�,,wn".^i�.��eF	BɉT��Qr�&�r�+0�+�V�b�LqY9��1	���Fc�9Y
���N��$V@�_Yq��y֘ŷ
A��o5������B�ϖ���]��3CR@5���>_��u ��I�:=]��H���h0��U�6l~�;D|��h���g�·���>�!�
���6�;~d,rЇ1h�<��qy_���.N�ܑ |O��Ca�Z����~y�H�3$>��Q�fZ(U_~��A&���Mg����(w�����X]��ol��B�0���+����0]5%�"|�K�1(`V�q�j�N��.�����]:�:�5�oPm�����{O3n��?R��dm|B���[����]m��݋C�ɿ	���^llp�s��h�:��$׭�4s�^�C��PB�A��6���]	��e�����9�!�P<y��!�˓�Ci�}'�Xq��!�z Qu���{��;(�,m��tl0W��A@67�HBI��9���*�a!�<7���x��Z�D �'�Qz�xf����-C���)Qo�.)���vN=��A�zM���g���?��(W�y�t�䦾�^짨�@O��e��K&caH��"'w3�����7��w/g�b�C�܆��ČLČ	�7U*����tͨr��%��;�-c�"Ö������b뚆f�D/6��վДCx�61�8l�1:Sr!��/�1��D�d6��?{K�N�21�]����o:R�Y�x���p�bP�p�O�;���0�����w$S�	i���